`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.11.2025 21:39:35
// Design Name: 
// Module Name: Mux_4x1_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mux_4x1_tb(
    );
     reg S1, S0, I0, I1, I2, I3;
    wire y;

    Mux_4x1 dut (S1, S0, I0, I1, I2, I3, y);

  initial begin
    S1=0; S0=0; I0=0; I1=0; I2=0; I3=0; #10;
    S1=0; S0=0; I0=0; I1=0; I2=0; I3=1; #10;
    S1=0; S0=0; I0=0; I1=0; I2=1; I3=0; #10;
    S1=0; S0=0; I0=0; I1=0; I2=1; I3=1; #10;
    S1=0; S0=0; I0=0; I1=1; I2=0; I3=0; #10;
    S1=0; S0=0; I0=0; I1=1; I2=0; I3=1; #10;
    S1=0; S0=0; I0=0; I1=1; I2=1; I3=0; #10;
    S1=0; S0=0; I0=0; I1=1; I2=1; I3=1; #10;
    S1=0; S0=0; I0=1; I1=0; I2=0; I3=0; #10;
    S1=0; S0=0; I0=1; I1=0; I2=0; I3=1; #10;
    S1=0; S0=0; I0=1; I1=0; I2=1; I3=0; #10;
    S1=0; S0=0; I0=1; I1=0; I2=1; I3=1; #10;
    S1=0; S0=0; I0=1; I1=1; I2=0; I3=0; #10;
    S1=0; S0=0; I0=1; I1=1; I2=0; I3=1; #10;
    S1=0; S0=0; I0=1; I1=1; I2=1; I3=0; #10;
    S1=0; S0=0; I0=1; I1=1; I2=1; I3=1; #10;
    S1=0; S0=1; I0=0; I1=0; I2=0; I3=0; #10;
    S1=0; S0=1; I0=0; I1=0; I2=0; I3=1; #10;
    S1=0; S0=1; I0=0; I1=0; I2=1; I3=0; #10;
    S1=0; S0=1; I0=0; I1=0; I2=1; I3=1; #10;
    S1=0; S0=1; I0=0; I1=1; I2=0; I3=0; #10;
    S1=0; S0=1; I0=0; I1=1; I2=0; I3=1; #10;
    S1=0; S0=1; I0=0; I1=1; I2=1; I3=0; #10;
    S1=0; S0=1; I0=0; I1=1; I2=1; I3=1; #10;
    S1=0; S0=1; I0=1; I1=0; I2=0; I3=0; #10;
    S1=0; S0=1; I0=1; I1=0; I2=0; I3=1; #10;
    S1=0; S0=1; I0=1; I1=0; I2=1; I3=0; #10;
    S1=0; S0=1; I0=1; I1=0; I2=1; I3=1; #10;
    S1=0; S0=1; I0=1; I1=1; I2=0; I3=0; #10;
    S1=0; S0=1; I0=1; I1=1; I2=0; I3=1; #10;
    S1=0; S0=1; I0=1; I1=1; I2=1; I3=0; #10;
    S1=0; S0=1; I0=1; I1=1; I2=1; I3=1; #10;
    S1=1; S0=0; I0=0; I1=0; I2=0; I3=0; #10;
    S1=1; S0=0; I0=0; I1=0; I2=0; I3=1; #10;
    S1=1; S0=0; I0=0; I1=0; I2=1; I3=0; #10;
    S1=1; S0=0; I0=0; I1=0; I2=1; I3=1; #10;
    S1=1; S0=0; I0=0; I1=1; I2=0; I3=0; #10;
    S1=1; S0=0; I0=0; I1=1; I2=0; I3=1; #10;
    S1=1; S0=0; I0=0; I1=1; I2=1; I3=0; #10;
    S1=1; S0=0; I0=0; I1=1; I2=1; I3=1; #10;
    S1=1; S0=0; I0=1; I1=0; I2=0; I3=0; #10;
    S1=1; S0=0; I0=1; I1=0; I2=0; I3=1; #10;
    S1=1; S0=0; I0=1; I1=0; I2=1; I3=0; #10;
    S1=1; S0=0; I0=1; I1=0; I2=1; I3=1; #10;
    S1=1; S0=0; I0=1; I1=1; I2=0; I3=0; #10;
    S1=1; S0=0; I0=1; I1=1; I2=0; I3=1; #10;
    S1=1; S0=0; I0=1; I1=1; I2=1; I3=0; #10;
    S1=1; S0=0; I0=1; I1=1; I2=1; I3=1; #10;
    S1=1; S0=1; I0=0; I1=0; I2=0; I3=0; #10;
    S1=1; S0=1; I0=0; I1=0; I2=0; I3=1; #10;
    S1=1; S0=1; I0=0; I1=0; I2=1; I3=0; #10;
    S1=1; S0=1; I0=0; I1=0; I2=1; I3=1; #10;
    S1=1; S0=1; I0=0; I1=1; I2=0; I3=0; #10;
    S1=1; S0=1; I0=0; I1=1; I2=0; I3=1; #10;
    S1=1; S0=1; I0=0; I1=1; I2=1; I3=0; #10;
    S1=1; S0=1; I0=0; I1=1; I2=1; I3=1; #10;
    S1=1; S0=1; I0=1; I1=0; I2=0; I3=0; #10;
    S1=1; S0=1; I0=1; I1=0; I2=0; I3=1; #10;
    S1=1; S0=1; I0=1; I1=0; I2=1; I3=0; #10;
    S1=1; S0=1; I0=1; I1=0; I2=1; I3=1; #10;
    S1=1; S0=1; I0=1; I1=1; I2=0; I3=0; #10;
    S1=1; S0=1; I0=1; I1=1; I2=0; I3=1; #10;
    S1=1; S0=1; I0=1; I1=1; I2=1; I3=0; #10;
    S1=1; S0=1; I0=1; I1=1; I2=1; I3=1; #10;
    $finish;
  end
endmodule
